module month_day(
		 input [3:0]  lsd,
		 input [3:0]  msd,
		 input [7:0]  count,
		 input 	      leap_year,
		 output [4:0] day,
		 output [3:0] month
		 );

   reg [4:0] 		      day_tmp;
   reg [3:0] 		      month_tmp;
   
   

   always @(lsd)
     begin
	
	if(count >= 91 + leap_year)
	  begin
	     month_tmp <= 4;
	     day_tmp <= count - (90 + leap_year);
	  end
	
	else if(count >= (60 + leap_year))
	  begin
	     month_tmp <= 3;
	     day_tmp <= count - (59 + leap_year);
	  end
	
	else if(count >= 32)
	  begin
	     month_tmp <= 2;
	     day_tmp <= count - 31;
	  end
	
	else
	  begin
	     month_tmp <= 1;
	     day_tmp <= count;
	  end
	
     end

   assign month = month_tmp;
   assign day = day_tmp;
   
   
endmodule // month_day


   
